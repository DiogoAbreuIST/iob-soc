assign gpio_input = 2000;
