assign gpio_input = 2022;
