assign gpio_input = 10;
assign DATA_IN = 406840;
