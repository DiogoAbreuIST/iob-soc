assign gpio_input = 10;
